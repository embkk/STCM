class Transaction;
  logic[15:0] data;
  logic[3:0] len;
endclass
package testbench_pkg;
  `include "transaction_tb.sv"
  `include "driver_tb.sv"
  `include "monitor_tb.sv"
    `include "scoreboard_tb.sv"
  `include "generator_tb.sv"
  `include "environment_tb.sv"
endpackage

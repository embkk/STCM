module serializer_tb #(
  parameters
) (
  input  logic  clk_i,
  input  logic  rst_i,
  output logic  tb_finished_o,
  output logic  tb_failed_o
);
  
endmodule
class Scoreboard;
task main();
endtask
endclass